--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package partido is
	constant NumeroPartidos : integer := 10 ;
	constant frecFPGA : integer := 50000000 ;
end partido ;

package body partido is
end partido ;
